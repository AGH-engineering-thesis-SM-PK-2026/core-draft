`define N_th_WORD_BEGIN(N)  (N*32)
`define N_th_STRB_BEGIN(N)  (N*4)

`define N_th_WORD_END(N)  (N*32 + 31)
`define N_th_STRB_END(N)  (N*4 + 3)