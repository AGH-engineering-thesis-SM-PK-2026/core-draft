`timescale 1ns / 1ps

// VGA terminal controller
// The terminal and CPU run in different clock domains, and it is necessary to
// cross clock domains safely. The module also converts ASCII to font glyphs'
// indices. The modules stores the current position of the virtual cursor,
// under which new characters will appear. The cursor can also be controlled
// by the user.
// The user can write to 4 locations:
// - WRITE1 (00) - write a character under the cursor
// - WRITEX (01) - change X position of cursor
// - WRITEY (10) - change Y position of cursor
// - WRITEA (11) - write attribute to the character under the cursor (not used)
// Szymon Miękina - 03.12.2025

module termctl (
    input wire          n_rst,
    input wire          cpuclk,     // CPU side clock signal
    input wire          vgaclk,     // VGA side clock signal
    input wire [1:0]    dstin,      // location write destination
    input wire [7:0]    datain,     // location write data
    input wire          trig,       // write trigger
    output reg          busy,       // controller busy writing to framebuffer
    output reg [6:0]    xwrite,     // write x component
    output reg [4:0]    ywrite,     // write y component
    input wire          writeack,   // write acknowledged by framebuffer
    output reg          writereq,   // write request to framebuffer
    output wire [7:0]   charout     // char out to framebuffer
);

wire nonprint;
wire newline;

wire [5:0] fontout;

// convert ASCII to glyph index
asciitofont tofont (
    .charin(datain),
    .fontout(fontout),
    .nonprint(nonprint),
    .newline(newline)   
);

// 00 color
assign charout = {2'b00, fontout};

reg [3:0] wrstate;

`define WR_INIT 4'b0000
`define WR_WRITE1 4'b0100
`define WR_WRITEX 4'b0101
`define WR_WRITEY 4'b0110
`define WR_WRITEA 4'b0111
`define WR_WAIT1 4'b1000
`define WR_WAITE 4'b1001
`define WR_NEXT1 4'b1010
`define WR_FINISH 4'b1111

// internal signals
reg u_writereq;
// metastable reg. (1st stage of 2FF synch.)
reg m_writereq;
reg m_writeack;
// synchronized reg. (2nd stage of 2FF synch.)
reg s_writeack;
// also writereq

always @(posedge cpuclk) begin
    case (wrstate)
    `WR_INIT: begin
        busy <= 1'b0;
        if (trig) begin
            busy <= 1'b1;
            wrstate <= `WR_WRITE1;
            case (dstin)
            2'b00: wrstate <= `WR_WRITE1;
            2'b01: wrstate <= `WR_WRITEX;
            2'b10: wrstate <= `WR_WRITEY;
            2'b11: wrstate <= `WR_WRITEA;
            endcase
        end
    end
    `WR_WRITE1: begin
        // write one char
        if (!nonprint) u_writereq <= 1'b1;
        wrstate <= `WR_WAIT1;
    end
    `WR_WRITEX: begin
        // update x
        xwrite <= datain[6:0];
        wrstate <= `WR_WAITE;
    end
    `WR_WRITEY: begin
        // update y
        ywrite <= datain[4:0];
        wrstate <= `WR_WAITE;
    end
    `WR_WRITEA: begin
        // write attribute (not used for now)
        wrstate <= `WR_WAITE;
    end
    `WR_WAIT1: begin
        // wait for the framebuffer to finish the char write
        u_writereq <= 1'b0;
        if (!s_writeack) wrstate <= `WR_NEXT1;
    end
    `WR_WAITE: begin
        wrstate <= `WR_FINISH;
    end
    `WR_NEXT1: begin
        // advance cursor to the next column or line
        xwrite <= xwrite + 1'b1;
        if (newline || xwrite == 99) begin
            ywrite <= ywrite + 1'b1;
            xwrite <= 1'b0;
        end
        wrstate <= `WR_FINISH;
    end
    `WR_FINISH: begin
        wrstate <= `WR_INIT;
        if (trig) wrstate <= `WR_FINISH;
    end
    endcase
    
    if (!n_rst) begin
        wrstate <= `WR_INIT;
        xwrite <= 1'b0;
        ywrite <= 1'b0;
    end
end


always @(posedge vgaclk) begin
    // writereq synchronizer
    m_writereq <= u_writereq;
    writereq <= m_writereq;
    
    // writeack synchronizer
    m_writeack <= writeack;
    s_writeack <= m_writeack;
end

endmodule
