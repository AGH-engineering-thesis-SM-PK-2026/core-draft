`timescale 1ns / 1ps

module toplevel(
    input       GLOBAL_CLK_IN
);

endmodule